`timescale 1ns / 1ps
/** @file AXIToStream_orchestrator.sv
 * @brief orchestrator top module Axi to axistream translation
 * @details
 * todo
 */

module AXIToStream_orchestrator_Reg #(
    parameter DATA_WIDTH = 128,
    parameter ADDR_WIDTH = 64,
    parameter ID_WIDTH = 32,
    parameter BURST_LEN = 8,
    parameter LOCK_WIDTH = 2,
    parameter USER_WIDTH = 64,
    parameter DEST_WIDTH = 32,
    localparam TIMER_WIDTH=DATA_WIDTH-ADDR_WIDTH-ID_WIDTH-BURST_LEN-channels_bits,
    // how many channels this module supports
    parameter channels = 6,
    //the bit needed to represent this channels in binary
    localparam channels_bits = $clog2(channels),

    localparam NONE_ID = 0,
    localparam AR_ID = 1,
    localparam AW_ID = 2,
    localparam R_ID = 3,
    localparam W_ID = 4,
    localparam B_ID = 5
  
) (
    input  wire                    clk,
    input  wire                    resetn,
    // reset params
    input wire [channels-1:0] submodule_resets,
    
    // AXI Slave (input wire) interface, will AXIS a transaction
    input  wire [    ID_WIDTH-1:0] AXIS_awid,
    input  wire [  ADDR_WIDTH-1:0] AXIS_awaddr,
    input  wire [   BURST_LEN-1:0] AXIS_awlen,
    input  wire [             2:0] AXIS_awsize,
    input  wire [             1:0] AXIS_awburst,
    input  wire [  LOCK_WIDTH-1:0] AXIS_awlock,
    input  wire [             3:0] AXIS_awcache,
    input  wire [             2:0] AXIS_awprot,
    input  wire [             3:0] AXIS_awregion,
    input  wire [             3:0] AXIS_awqos,
    input  wire [  USER_WIDTH-1:0] AXIS_awuser,
    input  wire                    AXIS_awvalid,
    output wire                    AXIS_awready,
    input  wire [    ID_WIDTH-1:0] AXIS_wid,
    input  wire [  DATA_WIDTH-1:0] AXIS_wdata,
    input  wire [DATA_WIDTH/8-1:0] AXIS_wstrb,
    input  wire                    AXIS_wlast,
    input  wire [  USER_WIDTH-1:0] AXIS_wuser,
    input  wire                    AXIS_wvalid,
    output wire                    AXIS_wready,
    output wire [    ID_WIDTH-1:0] AXIS_bid,
    output wire [             1:0] AXIS_bresp,
    output wire [  USER_WIDTH-1:0] AXIS_buser,
    output wire                    AXIS_bvalid,
    input  wire                    AXIS_bready,
    input  wire [    ID_WIDTH-1:0] AXIS_arid,
    input  wire [  ADDR_WIDTH-1:0] AXIS_araddr,
    input  wire [   BURST_LEN-1:0] AXIS_arlen,
    input  wire [             2:0] AXIS_arsize,
    input  wire [             1:0] AXIS_arburst,
    input  wire [  LOCK_WIDTH-1:0] AXIS_arlock,
    input  wire [             3:0] AXIS_arcache,
    input  wire [             2:0] AXIS_arprot,
    input  wire [             3:0] AXIS_arregion,
    input  wire [             3:0] AXIS_arqos,
    input  wire [  USER_WIDTH-1:0] AXIS_aruser,
    input  wire                    AXIS_arvalid,
    output wire                    AXIS_arready,
    output wire [    ID_WIDTH-1:0] AXIS_rid,
    output wire [  DATA_WIDTH-1:0] AXIS_rdata,
    output wire [             1:0] AXIS_rresp,
    output wire                    AXIS_rlast,
    output wire [  USER_WIDTH-1:0] AXIS_ruser,
    output wire                    AXIS_rvalid,
    input  wire                    AXIS_rready,
    // AXI master (output wire) Interface, will AXIM the AXISed transaction to destination
    output wire [    ID_WIDTH-1:0] AXIM_awid,
    output wire [  ADDR_WIDTH-1:0] AXIM_awaddr,
    output wire [   BURST_LEN-1:0] AXIM_awlen,
    output wire [             2:0] AXIM_awsize,
    output wire [             1:0] AXIM_awburst,
    output wire [  LOCK_WIDTH-1:0] AXIM_awlock,
    output wire [             3:0] AXIM_awcache,
    output wire [             2:0] AXIM_awprot,
    output wire [             3:0] AXIM_awregion,
    output wire [             3:0] AXIM_awqos,
    output wire [  USER_WIDTH-1:0] AXIM_awuser,
    output wire                    AXIM_awvalid,
    input  wire                    AXIM_awready,
    output wire [    ID_WIDTH-1:0] AXIM_wid,
    output wire [  DATA_WIDTH-1:0] AXIM_wdata,
    output wire [DATA_WIDTH/8-1:0] AXIM_wstrb,
    output wire                    AXIM_wlast,
    output wire [  USER_WIDTH-1:0] AXIM_wuser,
    output wire                    AXIM_wvalid,
    input  wire                    AXIM_wready,
    input  wire [    ID_WIDTH-1:0] AXIM_bid,
    input  wire [             1:0] AXIM_bresp,
    input  wire [  USER_WIDTH-1:0] AXIM_buser,
    input  wire                    AXIM_bvalid,
    output wire                    AXIM_bready,
    output wire [    ID_WIDTH-1:0] AXIM_arid,
    output wire [  ADDR_WIDTH-1:0] AXIM_araddr,
    output wire [   BURST_LEN-1:0] AXIM_arlen,
    output wire [             2:0] AXIM_arsize,
    output wire [             1:0] AXIM_arburst,
    output wire [  LOCK_WIDTH-1:0] AXIM_arlock,
    output wire [             3:0] AXIM_arcache,
    output wire [             2:0] AXIM_arprot,
    output wire [             3:0] AXIM_arregion,
    output wire [             3:0] AXIM_arqos,
    output wire [  USER_WIDTH-1:0] AXIM_aruser,
    output wire                    AXIM_arvalid,
    input  wire                    AXIM_arready,
    input  wire [    ID_WIDTH-1:0] AXIM_rid,
    input  wire [  DATA_WIDTH-1:0] AXIM_rdata,
    input  wire [             1:0] AXIM_rresp,
    input  wire                    AXIM_rlast,
    input  wire [  USER_WIDTH-1:0] AXIM_ruser,
    input  wire                    AXIM_rvalid,
    output wire                    AXIM_rready,
    // AXI stream Master (stream output wire) interface
    output wire [    ID_WIDTH-1:0] stream_tid,
    output wire [  DEST_WIDTH-1:0] stream_tdest,
    output reg [  DATA_WIDTH-1:0] stream_tdata,
    output wire [DATA_WIDTH/8-1:0] stream_tstrb,
    output wire [DATA_WIDTH/8-1:0] stream_tkeep,
    output reg                    stream_tlast,
    output wire [  USER_WIDTH-1:0] stream_tuser,
    output reg                    stream_tvalid,
    input  wire                    stream_tready

);
  //Submodules instantiation
  AXIToStream_Ax #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(ADDR_WIDTH),
      .ID_WIDTH(ID_WIDTH),
      .BURST_LEN(BURST_LEN),
      .LOCK_WIDTH(LOCK_WIDTH),
      .USER_WIDTH(USER_WIDTH),
      .STREAM_TYPE_WIDTH(channels_bits),
      .STREAM_TYPE(AR_ID),
      .TIMER_WIDTH(TIMER_WIDTH)
  ) AR (
      .clk(clk),
      .resetn(resets[AR_ID]),
      .ready(Orchestrator_ready[AR_ID]),
      .valid(submodule_valid[AR_ID]),
      .data(submodule_data[AR_ID]),
      .in_progress(submodule_in_progress[AR_ID]),
      .last(submodule_last[AR_ID]),
      .submodule_transaction_length(submodule_transaction_length[AR_ID]),
      .timestamp(timestamp),

      //subordinate
      .AXIS_axid(AXIS_arid),
      .AXIS_axaddr(AXIS_araddr),
      .AXIS_axlen(AXIS_arlen),
      .AXIS_axsize(AXIS_arsize),
      .AXIS_axburst(AXIS_arburst),
      .AXIS_axlock(AXIS_arlock),
      .AXIS_axcache(AXIS_arcache),
      .AXIS_axprot(AXIS_arprot),
      .AXIS_axregion(AXIS_arregion),
      .AXIS_axqos(AXIS_arqos),
      .AXIS_axuser(AXIS_aruser),
      .AXIS_axready(AXIS_arready),
      .AXIS_axvalid(AXIS_arvalid),

      //manager
      .AXIM_axid(AXIM_arid),
      .AXIM_axaddr(AXIM_araddr),
      .AXIM_axlen(AXIM_arlen),
      .AXIM_axsize(AXIM_arsize),
      .AXIM_axburst(AXIM_arburst),
      .AXIM_axlock(AXIM_arlock),
      .AXIM_axcache(AXIM_arcache),
      .AXIM_axprot(AXIM_arprot),
      .AXIM_axregion(AXIM_arregion),
      .AXIM_axqos(AXIM_arqos),
      .AXIM_axuser(AXIM_aruser),
      .AXIM_axready(AXIM_arready),
      .AXIM_axvalid(AXIM_arvalid)
  );

  AXIToStream_Ax #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(ADDR_WIDTH),
      .ID_WIDTH(ID_WIDTH),
      .BURST_LEN(BURST_LEN),
      .LOCK_WIDTH(LOCK_WIDTH),
      .USER_WIDTH(USER_WIDTH),
      .STREAM_TYPE_WIDTH(channels_bits),
      .STREAM_TYPE(AW_ID),
      .TIMER_WIDTH(TIMER_WIDTH)
  ) AW (
      .clk(clk),
      .resetn(resets[AW_ID]),
      .ready(Orchestrator_ready[AW_ID]),
      .valid(submodule_valid[AW_ID]),
      .data(submodule_data[AW_ID]),
      .in_progress(submodule_in_progress[AW_ID]),
      .last(submodule_last[AW_ID]),
      .submodule_transaction_length(submodule_transaction_length[AW_ID]),
      .timestamp(timestamp),

      //subordinate
      .AXIS_axid(AXIS_awid),
      .AXIS_axaddr(AXIS_awaddr),
      .AXIS_axlen(AXIS_awlen),
      .AXIS_axsize(AXIS_awsize),
      .AXIS_axburst(AXIS_awburst),
      .AXIS_axlock(AXIS_awlock),
      .AXIS_axcache(AXIS_awcache),
      .AXIS_axprot(AXIS_awprot),
      .AXIS_axregion(AXIS_awregion),
      .AXIS_axqos(AXIS_awqos),
      .AXIS_axuser(AXIS_awuser),
      .AXIS_axready(AXIS_awready),
      .AXIS_axvalid(AXIS_awvalid),

      //manager
      .AXIM_axid(AXIM_awid),
      .AXIM_axaddr(AXIM_awaddr),
      .AXIM_axlen(AXIM_awlen),
      .AXIM_axsize(AXIM_awsize),
      .AXIM_axburst(AXIM_awburst),
      .AXIM_axlock(AXIM_awlock),
      .AXIM_axcache(AXIM_awcache),
      .AXIM_axprot(AXIM_awprot),
      .AXIM_axregion(AXIM_awregion),
      .AXIM_axqos(AXIM_awqos),
      .AXIM_axuser(AXIM_awuser),
      .AXIM_axready(AXIM_awready),
      .AXIM_axvalid(AXIM_awvalid)
  );

  AXIToStream_B #(
      .DATA_WIDTH(DATA_WIDTH),
      .ID_WIDTH(ID_WIDTH),
      .USER_WIDTH(USER_WIDTH),
      .STREAM_TYPE_WIDTH(channels_bits),
      .STREAM_TYPE(B_ID)
  ) B (
      .clk(clk),
      .resetn(resets[B_ID]),
      .ready(Orchestrator_ready[B_ID]),
      .valid(submodule_valid[B_ID]),
      .data(submodule_data[B_ID]),
      .in_progress(submodule_in_progress[B_ID]),
      .last(submodule_last[B_ID]),
      .submodule_transaction_length(submodule_transaction_length[B_ID]),

      // AXI master (output wire) Interface, will forward the AXIS transaction to destination
      .AXIM_bid(AXIM_bid),
      .AXIM_bresp(AXIM_bresp),
      .AXIM_buser(AXIM_buser),
      .AXIM_bvalid(AXIM_bvalid),
      .AXIM_bready(AXIM_bready),
      // AXI Slave (input wire) interface
      .AXIS_bid(AXIS_bid),
      .AXIS_bresp(AXIS_bresp),
      .AXIS_buser(AXIS_buser),
      .AXIS_bvalid(AXIS_bvalid),
      .AXIS_bready(AXIS_bready)
  );

  Dummy_AXIToStream_R # (
      .DATA_WIDTH(DATA_WIDTH),
      .ID_WIDTH  (ID_WIDTH),
      .USER_WIDTH(USER_WIDTH)
      //.STREAM_TYPE_WIDTH(channels_bits),
      //.STREAM_TYPE(R_ID)
  ) R (
      .clk(clk),
      .resetn(resets[R_ID]),
      .ready(Orchestrator_ready[R_ID]),
      .valid(submodule_valid[R_ID]),
      .data(submodule_data[R_ID]),
      .in_progress(submodule_in_progress[R_ID]),
      .last(submodule_last[R_ID]),
      .submodule_transaction_length(submodule_transaction_length[R_ID]),
      // AXI master (output wire) Interface, will forward the AXIS transaction to destination
      .AXIM_rid(AXIM_rid),
      .AXIM_rdata(AXIM_rdata),
      .AXIM_rresp(AXIM_rresp),
      .AXIM_rlast(AXIM_rlast),
      .AXIM_ruser(AXIM_ruser),
      .AXIM_rvalid(AXIM_rvalid),
      .AXIM_rready(AXIM_rready),
      // AXI Slave (input wire) interface
      .AXIS_rid(AXIS_rid),
      .AXIS_rdata(AXIS_rdata),
      .AXIS_rresp(AXIS_rresp),
      .AXIS_rlast(AXIS_rlast),
      .AXIS_ruser(AXIS_ruser),
      .AXIS_rvalid(AXIS_rvalid),
      .AXIS_rready(AXIS_rready)
  );

  

  Dummy_AXIToStream_W #(
      .DATA_WIDTH(DATA_WIDTH),
      .ID_WIDTH  (ID_WIDTH),
      .USER_WIDTH(USER_WIDTH)
      //.STREAM_TYPE_WIDTH(channels_bits),
      //.STREAM_TYPE(W_ID),
      //.BURST_SIZE(BURST_LEN)
  ) W (
      .clk(clk),
      .resetn(resets[W_ID]),
      .ready(Orchestrator_ready[W_ID]),
      .valid(submodule_valid[W_ID]),
      .data(submodule_data[W_ID]),
      .in_progress(submodule_in_progress[W_ID]),
      .last(submodule_last[W_ID]),
      .submodule_transaction_length(submodule_transaction_length[W_ID]),
      // AXI master (output wire) Interface, will forward the AXIS transaction to destination
      .AXIM_wid(AXIM_wid),
      .AXIM_wdata(AXIM_wdata),
      .AXIM_wstrb(AXIM_wstrb),
      .AXIM_wlast(AXIM_wlast),
      .AXIM_wuser(AXIM_wuser),
      .AXIM_wvalid(AXIM_wvalid),
      .AXIM_wready(AXIM_wready),
      // AXI Slave (input wire) interface
      .AXIS_wid(AXIS_wid),
      .AXIS_wdata(AXIS_wdata),
      .AXIS_wstrb(AXIS_wstrb),
      .AXIS_wlast(AXIS_wlast),
      .AXIS_wuser(AXIS_wuser),
      .AXIS_wvalid(AXIS_wvalid),
      .AXIS_wready(AXIS_wready)
  );
  reg [channels_bits:0] State;//interpret this as last
  reg [TIMER_WIDTH-1:0] timestamp;

  //AXI stream wirings
  assign stream_tid   = 0;
  assign stream_tdest = 0;
  assign stream_tstrb = 0;
  assign stream_tkeep = {DATA_WIDTH / 8{1'b1}};
  assign stream_tuser = 0;

  wire[channels-1:0][channels-1:0] encodings;

//all the unused channels have their ready,last,valid and in_progress to 0


  ///send reset to individual submodules (and keep unwanted submodules in reset)
  wire [channels-1:0] resets;
  assign resets[AR_ID] = resetn && submodule_resets[AR_ID];
  assign resets[AW_ID] = resetn && submodule_resets[AW_ID];
  assign resets[R_ID]  = resetn && submodule_resets[R_ID];
  assign resets[W_ID]  = resetn && submodule_resets[W_ID];
  assign resets[B_ID]  = resetn && submodule_resets[B_ID];

  /// how the top module signals a specific submodule that the transaction can proceed
  reg [channels-1:0] Orchestrator_ready;

  /// how the submodules will signal to the top module that they have valid data
  /// (after having detected a handshake between the two original axi
  /// interfaces), or a multi-clock cycle transaction is still in progress (e.g.
  /// R/w).
  wire [channels-1:0] submodule_valid, submodule_in_progress, submodule_last;
  //the next to have the data
  wire [channels-1:0][DATA_WIDTH-1:0] submodule_data;
  wire [channels-1:0][5:0]submodule_transaction_length;

  ///to implement round robin we need a register that will cycle between all the
  ///possible channels (when they are valid)
  // this register will hold the id of the last channel that has transmitted
  // data
  //reg [channels_bits-1:0] last_index;
  
  genvar k;
  generate
   for (k = 0; k < channels; k++) begin
      //Make first encoding all 0 for NONE state
      if(k>0)begin
        assign encodings[k] = {{channels{1'b0}} | {1'b1}}<<k;
      end
      else begin
        assign encodings[k] = {channels{1'b0}};
        
      end
   end
   endgenerate

        assign submodule_data[0]=0;
        assign submodule_in_progress[0]=0;
        assign submodule_last[0]=0;
        assign submodule_valid[0]=0;
        assign resets[0]=1;
        assign submodule_transaction_length[0]=0;
        //assign submodule_resets[0]=0;

  reg [5:0] transaction_length;
 
  //stateChanger!
  integer i=0;
//  always @(posedge clk) begin
//    if (!resetn) begin
//    //last_index<=0;
//    State<=0;
//    timestamp<=0;
//    end
//    else begin
//      //if the state that we were in last is still performing a transaction and/or downstream is not ready then do not change states 
//      if (~submodule_in_progress[State] & transaction_length==0)  begin
//        //check if any submodules have data pending
//        if(|submodule_valid)begin
//          //change state to the next submodule that has valid data waiting to be sent
//          for (i = 1; i <=channels; i++) begin 
//            //explicitly check to wrap around when checking who is the first valid submodule
//            if (submodule_valid[(State+i>channels) ? (State+i-channels):(State+i)])begin
//               //change the state when the first valid submodule is found
//               State<=(State+i>channels) ? (State+i-channels):(State+i);
//               break;
//            end
//          end
//        end
//        //if no submodule ready, then switch to the NONE State
//        // else begin
//        //   State<=0;
//        // end
//      end
//      //state is in progress. update something 
//      else begin
//        State<=State;
//      end
//      timestamp<=timestamp+1;
//    end

//  end
  
  reg [channels_bits:0] NextState;
  
  always @(posedge clk) begin
    if (!resetn) begin
    //last_index<=0;
    State<=0;
    timestamp<=0;
    
    end
    else begin
      State<=NextState;
      timestamp<=timestamp+1;
    end

  end
  
  always @* begin 
  if (!resetn) begin
  NextState<=0;
  end
  if (~submodule_in_progress[State] & transaction_length==0)  begin
        //check if any submodules have data pending
        if(|submodule_valid)begin
          //change state to the next submodule that has valid data waiting to be sent
          for (i = 1; i <=channels; i++) begin 
            //explicitly check to wrap around when checking who is the first valid submodule
            if (submodule_valid[(State+i>channels) ? (State+i-channels):(State+i)])begin
               //change the state when the first valid submodule is found
               NextState<=(State+i>channels) ? (State+i-channels):(State+i);
               break;
            end
          end
        end
  end
  end
  
  reg started;
  //DATAMOVER!
  int j;
  //this block will handle AXISTREAM and Submodule Orchestration
  always @(posedge clk) begin
    if(!resetn)begin
      Orchestrator_ready<=encodings[0];
      stream_tdata<=0;
      stream_tlast<=0;
      stream_tvalid<=0;
      transaction_length<=0;
      started<=0;
    end
    else begin
      if(State!=0 & stream_tready)begin
        if(transaction_length>=1 & started)begin
          //start the transaction
          Orchestrator_ready<=encodings[State];                             
          stream_tdata<=submodule_data[State];
          stream_tlast<=submodule_last[State];
          stream_tvalid<=1;
          transaction_length<=transaction_length-1;
        end
        else if (transaction_length==0 & started) begin
          Orchestrator_ready<=encodings[0];
          stream_tdata<=0;
          stream_tlast<=0;
          stream_tvalid<=0;
          transaction_length<=0;
          started<=0;
        end
        else if (!started & submodule_valid[State])begin
          //grab the length
          transaction_length<=submodule_transaction_length[State];
          started<=1;
        end
        
      end
      else begin
        Orchestrator_ready<=encodings[0];
        stream_tdata<=0;
        stream_tlast<=0;
        stream_tvalid<=0;
        transaction_length<=0;
        started<=0;
      end
    end
  end

endmodule