`timescale 1ns / 1ps
/** @file AXIToStream.sv
 * @brief Snoop AXI4 transaction and send a copy of their data from the
 *  AXIStream port.
 * @author Mattia Nicolella
 */

/** @brief Snoop AXI4 transaction and send a copy of their data from the
 *  AXIStream port.
 * @details This module acts as a passtrough between an AXI4 master/slave,
 * while creating an equivalent transaction from the AXIStream master.
 *
 * *NOTE:* This module introduces a ~3 clock delay in each AXI4 transaction.
 */
module AXIToStream #(
    parameter DATA_WIDTH = 128,
    parameter ADDR_WIDTH = 64,
    parameter ID_WIDTH = 32,
    parameter BURST_LEN = 8,
    parameter LOCK_WIDTH = 2,
    parameter USER_WIDTH = 64,
    parameter DEST_WIDTH = 32,
    parameter STREAM_TYPE_WIDTH = 3,
    localparam STREAM_DATA_WIDTH = DATA_WIDTH + STREAM_TYPE_WIDTH + ADDR_WIDTH + (DATA_WIDTH / 8)
) (
    input  wire                    clk,
    input  wire                    resetn,
    // AXI Slave (input wire) interface, will snoop a transaction
    input  wire [    ID_WIDTH-1:0] snoop_awid,
    input  wire [  ADDR_WIDTH-1:0] snoop_awaddr,
    input  wire [   BURST_LEN-1:0] snoop_awlen,
    input  wire [             2:0] snoop_awsize,
    input  wire [             1:0] snoop_awburst,
    input  wire [  LOCK_WIDTH-1:0] snoop_awlock,
    input  wire [             3:0] snoop_awcache,
    input  wire [             2:0] snoop_awprot,
    input  wire [             3:0] snoop_awregion,
    input  wire [             3:0] snoop_awqos,
    input  wire [  USER_WIDTH-1:0] snoop_awuser,
    input  wire                    snoop_awvalid,
    output wire                    snoop_awready,
    input  wire [    ID_WIDTH-1:0] snoop_wid,
    input  wire [  DATA_WIDTH-1:0] snoop_wdata,
    input  wire [DATA_WIDTH/8-1:0] snoop_wstrb,
    input  wire                    snoop_wlast,
    input  wire [  USER_WIDTH-1:0] snoop_wuser,
    input  wire                    snoop_wvalid,
    output wire                    snoop_wready,
    output wire [    ID_WIDTH-1:0] snoop_bid,
    output wire [             1:0] snoop_bresp,
    output wire [  USER_WIDTH-1:0] snoop_buser,
    output wire                    snoop_bvalid,
    input  wire                    snoop_bready,
    input  wire [    ID_WIDTH-1:0] snoop_arid,
    input  wire [  ADDR_WIDTH-1:0] snoop_araddr,
    input  wire [   BURST_LEN-1:0] snoop_arlen,
    input  wire [             2:0] snoop_arsize,
    input  wire [             1:0] snoop_arburst,
    input  wire [  LOCK_WIDTH-1:0] snoop_arlock,
    input  wire [             3:0] snoop_arcache,
    input  wire [             2:0] snoop_arprot,
    input  wire [             3:0] snoop_arregion,
    input  wire [             3:0] snoop_arqos,
    input  wire [  USER_WIDTH-1:0] snoop_aruser,
    input  wire                    snoop_arvalid,
    output wire                    snoop_arready,
    output wire [    ID_WIDTH-1:0] snoop_rid,
    output wire [  DATA_WIDTH-1:0] snoop_rdata,
    output wire [             1:0] snoop_rresp,
    output wire                    snoop_rlast,
    output wire [  USER_WIDTH-1:0] snoop_ruser,
    output wire                    snoop_rvalid,
    input  wire                    snoop_rready,
    // AXI master (output wire) Interface, will forward the snooped transaction to destination
    output wire [    ID_WIDTH-1:0] forward_awid,
    output wire [  ADDR_WIDTH-1:0] forward_awaddr,
    output wire [   BURST_LEN-1:0] forward_awlen,
    output wire [             2:0] forward_awsize,
    output wire [             1:0] forward_awburst,
    output wire [  LOCK_WIDTH-1:0] forward_awlock,
    output wire [             3:0] forward_awcache,
    output wire [             2:0] forward_awprot,
    output wire [             3:0] forward_awregion,
    output wire [             3:0] forward_awqos,
    output wire [  USER_WIDTH-1:0] forward_awuser,
    output wire                    forward_awvalid,
    input  wire                    forward_awready,
    output wire [    ID_WIDTH-1:0] forward_wid,
    output wire [  DATA_WIDTH-1:0] forward_wdata,
    output wire [DATA_WIDTH/8-1:0] forward_wstrb,
    output wire                    forward_wlast,
    output wire [  USER_WIDTH-1:0] forward_wuser,
    output wire                    forward_wvalid,
    input  wire                    forward_wready,
    input  wire [    ID_WIDTH-1:0] forward_bid,
    input  wire [             1:0] forward_bresp,
    input  wire [  USER_WIDTH-1:0] forward_buser,
    input  wire                    forward_bvalid,
    output wire                    forward_bready,
    output wire [    ID_WIDTH-1:0] forward_arid,
    output wire [  ADDR_WIDTH-1:0] forward_araddr,
    output wire [   BURST_LEN-1:0] forward_arlen,
    output wire [             2:0] forward_arsize,
    output wire [             1:0] forward_arburst,
    output wire [  LOCK_WIDTH-1:0] forward_arlock,
    output wire [             3:0] forward_arcache,
    output wire [             2:0] forward_arprot,
    output wire [             3:0] forward_arregion,
    output wire [             3:0] forward_arqos,
    output wire [  USER_WIDTH-1:0] forward_aruser,
    output wire                    forward_arvalid,
    input  wire                    forward_arready,
    input  wire [    ID_WIDTH-1:0] forward_rid,
    input  wire [  DATA_WIDTH-1:0] forward_rdata,
    input  wire [             1:0] forward_rresp,
    input  wire                    forward_rlast,
    input  wire [  USER_WIDTH-1:0] forward_ruser,
    input  wire                    forward_rvalid,
    output wire                    forward_rready,
    // AXI stream Master (stream output wire) interface
    output wire [    ID_WIDTH-1:0] stream_tid,
    output wire [  DEST_WIDTH-1:0] stream_tdest,
    output wire [  DATA_WIDTH-1:0] stream_tdata,
    output wire [DATA_WIDTH/8-1:0] stream_tstrb,
    output wire [DATA_WIDTH/8-1:0] stream_tkeep,
    output wire                    stream_tlast,
    output wire [  USER_WIDTH-1:0] stream_tuser,
    output wire                    stream_tvalid,
    input  wire                    stream_tready,

    //debug pins
    output wire  DBG_can_forwardAR,
    output wire  DBG_can_forwardAW,
    output wire  DBG_can_forwardR,
    output wire  DBG_can_forwardW,
    output wire  DBG_can_forwardB
);

  /** The type of the ongoing stream (matches the AXI4 channels).
	 * *NOTE*: Each stream transaction is "tagged" with ::_stream_type so we need
	 * two bursts to send the read and write data. Additionally, the write data
	 * contains the original AXI4 strobe.
	 */
  enum reg [STREAM_TYPE_WIDTH-1:0] {
    NONE = 0,
    AR,
    R,
    AW,
    WSTRB,
    W,
    B
  } _stream_type;

  /** This register is used to make sure that we don´t starve neither read or write transactions,
   * by remembering which transaction was streamed during last contentions.
	 */
  enum reg [1:0] {
    NOC = 0,     //no conflict
    CAR,    // contention, do AR
    CAW    // contention, do AW
  } _address_rr;

  /** Data to be streamed in to the AXIStream slave.
   * In case of RDATA and WDATA streams we need to compose the metadata and
   * save the contents of the data line since we do not have any spare bits
   * in stream_tdata, so we use a tag team of two registers to send the output
   * save the one we will send next.
  */
  reg [DATA_WIDTH-1:0] _stream_data, _stream_data_next;

  /// Since we are deferring the data transaction we need to save its strobe to send them together
  reg [DATA_WIDTH/8-1:0] _stream_strobe;

  /**@brief keep track how how long is the burst,
   * reminder: burst len is defined as 1+Ax_LEN, and for R/W transaction
   */
  reg [BURST_LEN+1-1:0] _burst_len;


   //reg _data_sent
   //assign 


  /** To have meaningful transactions and not lose data we stall the AXI4 slave
	 * ready signal until the current AXIStream transaction has completed and
	 * the AXIStream is ready to process another transaction.
	 * We also ahve to enforce the AXI4 protocol dependencies for the different transactions
	 */
  /** We accept an AR transaction if:
	 * - stream module is ready (`stream_tready`)
	 * - we are not streaming already another transaction (`_stream_type==NONE`)
	 * - there is no conflict with a write transaction (`!snoop_arvalid`)
	 * - there was a conflict with a write transaction and we stalled the read transaction (`_address_rr == AW`)
	 */
  wire can_forwardAR;
  assign can_forwardAR = ~resetn || (stream_tready && _stream_type == NONE && (!snoop_awvalid || _address_rr != CAR));
  /** We accept an AW transaction if:
	 * - stream module is ready (`stream_tready`)
	 * - we are not streaming already another transaction (`_stream_type==NONE`)
	 * - there is no conflict with a write transaction (`!snoop_arvalid`)
	 * - there was a conflict with a write transaction and we stalled the read transaction (`_address_rr == AW`)
	 */
  wire can_forwardAW;
  assign can_forwardAW = ~resetn || (stream_tready && _stream_type == NONE && (!snoop_arvalid || _address_rr != CAW));
  ///For R/W  we depend on the completion of the previous AR/AW and there can be multiple R/W bursts in the same transaction
  wire can_forwardR, can_forwardW;
  assign can_forwardR = ~resetn || (stream_tready && (_stream_type == AR || _stream_type == R));
  assign can_forwardW = ~resetn || (stream_tready && _stream_type == WSTRB );
  /// For B transaction we only depend on the completion of the previous write transaction
  wire can_forwardB;
  assign can_forwardB = ~resetn || (stream_tready && _stream_type == W && _burst_len ==0);
  assign DBG_can_forwardAR = can_forwardAR;
  assign DBG_can_forwardR = can_forwardR;
  assign DBG_can_forwardAW = can_forwardAW;
  assign DBG_can_forwardW = can_forwardW;
  assign DBG_can_forwardB = can_forwardB;
  
  // connect the master to the slave port, so we can forward downstream the signals we received.
  assign forward_awid = snoop_awid;
  assign forward_awaddr = snoop_awaddr;
  assign forward_awlen = snoop_awlen;
  assign forward_awsize = snoop_awsize;
  assign forward_awburst = snoop_awburst;
  assign forward_awlock = snoop_awlock;
  assign forward_awcache = snoop_awcache;
  assign forward_awprot = snoop_awprot;
  assign forward_awregion = snoop_awregion;
  assign forward_awqos = snoop_awqos;
  assign forward_awuser = snoop_awuser;
  assign forward_awvalid = snoop_awvalid;
  assign snoop_awready = forward_awready;

  assign forward_wid = snoop_wid;
  assign forward_wdata = snoop_wdata;
  assign forward_wstrb = snoop_wstrb;
  assign forward_wlast = snoop_wlast;
  assign forward_wuser = snoop_wuser;
  assign forward_wvalid = snoop_wvalid;
  assign snoop_wready = forward_wready;

  assign snoop_bid = forward_bid;
  assign snoop_bresp = forward_bresp;
  assign snoop_buser = forward_buser;
  assign forward_bready = snoop_bready;
  assign snoop_bvalid = forward_bvalid;

  assign forward_arid = snoop_arid;
  assign forward_araddr = snoop_araddr;
  assign forward_arlen = snoop_arlen;
  assign forward_arsize = snoop_arsize;
  assign forward_arburst = snoop_arburst;
  assign forward_arlock = snoop_arlock;
  assign forward_arcache = snoop_arcache;
  assign forward_arprot = snoop_arprot;
  assign forward_arregion = snoop_arregion;
  assign forward_arqos = snoop_arqos;
  assign forward_aruser = snoop_aruser;
  assign forward_arvalid = snoop_arvalid && can_forwardAR;
  assign snoop_arready = forward_arready && can_forwardAR;

  assign snoop_rid = forward_rid;
  assign snoop_rdata = forward_rdata;
  assign snoop_rresp = forward_rresp;
  assign snoop_rlast = forward_rlast;
  assign snoop_ruser = forward_ruser;
  assign snoop_rvalid = forward_rvalid && can_forwardR;
  assign forward_rready = snoop_rready && can_forwardR;

  //state machine handling
  // we are using the valid and ready wires that take the streaming module state into account
  always @(posedge clk) begin
    if (~resetn) begin
      _stream_type <= NONE;
      _address_rr  <= NOC;
      _burst_len<=0;
      // Ax transaction
    end else if ((snoop_arvalid && forward_arready && can_forwardAR) || (snoop_awvalid && forward_awready && can_forwardAW)) begin
//        if((snoop_arvalid && forward_arready) && (snoop_awvalid && forward_awready) && _address_rr==NOC) //no conflict initially but then contention
//            _address_rr  <= (snoop_arvalid && forward_arready) ? CAR : CAW;//preference towards read going first
//        else begin
//            _address_rr <= NOC;
//        end
          _stream_type <= (snoop_arvalid && forward_arready) ? AR : AW;
          // arlen value + 1st burst transaction (manual specification) + metadata
          _burst_len   <= ((snoop_arvalid && forward_arready) ? snoop_arlen : snoop_awlen)+1+1;
          // R transaction
        end else if ((_stream_type==AR || _stream_type==R && can_forwardR) && ((snoop_rready && forward_rvalid)  || _burst_len == 1 )) begin
          _stream_type <= R;
          _address_rr  <= _address_rr;
          // we do not decrement the burst length if we are streaming AR
          _burst_len <= (_stream_type==AR)? _burst_len : _burst_len-1;
          // W transaction, here we grab the metadata and send it
        end 
//        else if (snoop_wready && forward_wvalid && can_forwardW && (_stream_type==AW || _stream_type ==W)) begin
//         _stream_type<=WSTRB;
//         _address_rr <=_address_rr;
//         _burst_len <= _burst_len;
//         // W transaction, send the actual data and prepare meteadata for next W burst
//         end 
//         else if (( snoop_wready && forward_wvalid && can_forwardW) || (_burst_len == 1 && can_forwardW)) begin
//         _stream_type <=W;
//         _address_rr <= _address_rr;
//         _burst_len <= _burst_len-1;      
//        end 
//        else if (snoop_bready && forward_bvalid && can_forwardB) begin
//          _stream_type <= B;
//          _burst_len   <= 0;
//          _address_rr  <= _address_rr;
//        end 
        else if (_burst_len == 0 && stream_tready && (_stream_type == R || _stream_type == B)) begin
          _stream_type <= (_stream_type == R || _stream_type == B) ? NONE : _stream_type;
          _burst_len   <= 0;
        end 
        else begin
          _stream_type <= _stream_type;
          _burst_len   <= _burst_len;
          _address_rr  <= _address_rr;
        end
  end


  //@bug: THIS HAS TO BE TOTALLY REWORKED ACCORDING TO THE STATE MACHINE ABOVE
	//build the stream data register
  always @(posedge clk) begin
    // reset
    if (~resetn) begin
        
      _stream_strobe <= 0;
      _stream_data <= 0;
      _stream_data_next <= 0;
      
    end
    // we are completing a single burst transaction, so we will go idle next clock
//    else if (((snoop_rready && _stream_type == R) || ( forward_wready && _stream_type == W)) && _burst_len==1) begin
      
//      _stream_data <= _stream_data_next;
//      _stream_data_next <= {DATA_WIDTH - 1{1'b0}};
//      _stream_strobe <= {DATA_WIDTH / 8{1'b1}};
//      // we are waiting for one interface
//    end
    //last element of R and W
    //questioning validity of below
    //barely makes it
    else if (_burst_len == 0 && stream_tready && (_stream_type == R || _stream_type == W)) begin
         _stream_data<=_stream_data_next;
         _stream_data_next<=0;
    end 
    /* transaction on the AR channel, pack the address with metadata and stream it
    *   stream what transaction is happening then pad with 0 then add the address
    *   burst lenght always has to be stated?
    */
    else if (snoop_arvalid && forward_arready && can_forwardAR) begin
      _stream_data <= {AR, {(DATA_WIDTH - STREAM_TYPE_WIDTH - ADDR_WIDTH) {1'b0}}, snoop_araddr};
      _stream_data_next <= {R, {(DATA_WIDTH - STREAM_TYPE_WIDTH) {1'b0}}};
      _stream_strobe <= {
        {(STREAM_TYPE_WIDTH + 7) / 8{1'b1}},
        {(DATA_WIDTH - STREAM_TYPE_WIDTH + 7 - ADDR_WIDTH) / 8{1'b0}},
        {ADDR_WIDTH / 8{1'b1}}
      };
      
    end 
    /* transaction on the AW channel, pack the address with metadata and stream it
    *   stream what transaction is happening then pad with 0 then add the address
    *
    */
    else if (snoop_awvalid && forward_awready && can_forwardAW) begin
      _stream_data <= {AW, {DATA_WIDTH - STREAM_TYPE_WIDTH - ADDR_WIDTH{1'b0}}, snoop_awaddr};
     
      _stream_strobe <= {
        {(STREAM_TYPE_WIDTH + 7) / 8{1'b1}},
        {(DATA_WIDTH - STREAM_TYPE_WIDTH + 7 - ADDR_WIDTH) / 8{1'b0}},
        {ADDR_WIDTH / 8{1'b1}}
      };
      
      // transaction on the B channel, pack resp with metadata and stream
    end 
    /* transaction on the B channel, pack the address with metadata and stream it
    *   stream what transaction is happening then pad with 0 then add the address
    *
    */
//    else if (snoop_bready && forward_bvalid && can_forwardB) begin
//      _stream_data <= {B, {DATA_WIDTH - STREAM_TYPE_WIDTH - 2{1'b0}}, snoop_bresp};
      
//      _stream_strobe <= {
//        {(STREAM_TYPE_WIDTH + 7) / 8{1'b1}},
//        {(DATA_WIDTH - STREAM_TYPE_WIDTH + 7 - 2) / 8{1'b0}},
//        8'b1
//      };
//      // 
//    end 
    /* 1st burst element of a transaction in the R channel, send the metadata created in the AR state and stored the data register
    * i.e. send metadata first, save the incoming data, then next clock cycle send the actual data
    *  NEEDS TO CHECK IF IT IS THE FIRST TIME GETTING R TRANSACTION
    */
    else if (snoop_rready &&  forward_rvalid && can_forwardR && _stream_type==AR) begin
     _stream_data <= _stream_data_next;
      _stream_data_next <= forward_rdata;
      _stream_strobe <= {
        {(STREAM_TYPE_WIDTH + 7) / 8{1'b1}}, {(DATA_WIDTH - STREAM_TYPE_WIDTH + 7) / 8{1'b0}}
      };
      // R transaction, from after sending the metadata
      // send the previous data burst and store the next
    end 
    else if (forward_rready &&  snoop_rvalid && can_forwardR && _stream_type==R) begin
      // the next state depends on forward_rlast
      
      _stream_data <= _stream_data_next;
      _stream_data_next <= forward_rdata;
      _stream_strobe <= {DATA_WIDTH{1'b1}};
      // last element of a burst transaction on the R channel
    end
//    //***something is supsicious about this conditional*** 
//    else if (forward_rready &&  snoop_rvalid && forward_rlast) begin
//      _stream_data <= _stream_data_next;
//      _stream_data_next <= {DATA_WIDTH - 1{1'b0}};
//      _stream_strobe <= {DATA_WIDTH / 8{1'b1}};
//      end
//      // Burst element of a transaction in the W channel, send the metadata and store the data
//    else if (forward_wready && snoop_wvalid && (_stream_type==AW ||_stream_type == W)) begin
   
//      _stream_data <= {W, {DATA_WIDTH - (DATA_WIDTH / 8) {1'b0}}, snoop_wstrb};
//      _stream_data_next <= snoop_wdata;
      
//      _stream_strobe <= {
//        {(STREAM_TYPE_WIDTH + 7) / 8{1'b1}},
//        {(DATA_WIDTH - STREAM_TYPE_WIDTH + 7 - DATA_WIDTH / 8) / 8{1'b0}},
//        {DATA_WIDTH / 8{1'b1}}
//      };
//      // W transaction, from after we sent the strobe
//      // send the previous data
//    end 
//    else if (can_forwardW) begin
//      // the next state depends on forward_rlast
      
//      _stream_data_next <=0; // only to avoid latching
//      _stream_data <= _stream_data_next;
//      _stream_strobe <= {DATA_WIDTH / 8{1'b1}};
//      // last element of a burst transaction on the W channel
//    end 
    else begin
      _stream_data <= _stream_data;
      _stream_data_next <= _stream_data_next;
      _stream_strobe <= _stream_strobe;
    end
  end

  // check wether the last piece of data was received
//  always @(posedge clk) begin
//    if (~resetn) begin
//      _stream_received <= 1;  // there's no data to send at reset
//    end else if (stream_tvalid && stream_tready) begin
//      _stream_received <= 1;
//    end else begin
//      _stream_received <= 0;
//    end
//  end


  // connect remaining AXI stream cables
  assign stream_tvalid = (can_forwardAR || can_forwardR) && _stream_type!=NONE;
  assign stream_tdata = _stream_data;
  assign stream_tstrb = _stream_strobe;
  assign stream_tkeep = {DATA_WIDTH / 8{1'b1}};
  assign stream_tlast = stream_tvalid && _burst_len==0;
  assign stream_tid = 0;
  assign stream_tdest = 0;
  assign stream_tuser = 0;
endmodule
