`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/14/2024 10:55:52 AM
// Design Name: 
// Module Name: AXIToStream_orchestrator_wrapper
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AXIToStream_orchestrator_wrapper#(
    parameter DATA_WIDTH = 128,
    parameter ADDR_WIDTH = 64,
    parameter ID_WIDTH = 32,
    parameter BURST_LEN = 8,
    parameter LOCK_WIDTH = 2,
    parameter USER_WIDTH = 64,
    parameter DEST_WIDTH = 32, 
    parameter CHANNELS = 6
)(
    input  wire                    clk,
    input  wire                    resetn,
    // AXI Slave (input wire) interface, will AXIS a transaction
    // input  wire                    RESETN_AR,
    // input  wire                    RESETN_AW,
    // input  wire                    RESETN_R,
    // input  wire                    RESETN_W,
    // input  wire                    RESETN_B,

    input wire [CHANNELS-1:0] submodule_resets,
         
    input  wire [    ID_WIDTH-1:0] AXIS_awid,
    input  wire [  ADDR_WIDTH-1:0] AXIS_awaddr,
    input  wire [   BURST_LEN-1:0] AXIS_awlen,
    input  wire [             2:0] AXIS_awsize,
    input  wire [             1:0] AXIS_awburst,
    input  wire [  LOCK_WIDTH-1:0] AXIS_awlock,
    input  wire [             3:0] AXIS_awcache,
    input  wire [             2:0] AXIS_awprot,
    input  wire [             3:0] AXIS_awregion,
    input  wire [             3:0] AXIS_awqos,
    input  wire [  USER_WIDTH-1:0] AXIS_awuser,
    input  wire                    AXIS_awvalid,
    output wire                    AXIS_awready,
    
    output wire [    ID_WIDTH-1:0] AXIM_awid,
    output wire [  ADDR_WIDTH-1:0] AXIM_awaddr,
    output wire [   BURST_LEN-1:0] AXIM_awlen,
    output wire [             2:0] AXIM_awsize,
    output wire [             1:0] AXIM_awburst,
    output wire [  LOCK_WIDTH-1:0] AXIM_awlock,
    output wire [             3:0] AXIM_awcache,
    output wire [             2:0] AXIM_awprot,
    output wire [             3:0] AXIM_awregion,
    output wire [             3:0] AXIM_awqos,
    output wire [  USER_WIDTH-1:0] AXIM_awuser,
    output wire                    AXIM_awvalid,
    input  wire                    AXIM_awready,
    
    input  wire [    ID_WIDTH-1:0] AXIS_wid,
    input  wire [  DATA_WIDTH-1:0] AXIS_wdata,
    input  wire [DATA_WIDTH/8-1:0] AXIS_wstrb,
    input  wire                    AXIS_wlast,
    input  wire [  USER_WIDTH-1:0] AXIS_wuser,
    input  wire                    AXIS_wvalid,
    output wire                    AXIS_wready,
    
    output wire [    ID_WIDTH-1:0] AXIM_wid,
    output wire [  DATA_WIDTH-1:0] AXIM_wdata,
    output wire [DATA_WIDTH/8-1:0] AXIM_wstrb,
    output wire                    AXIM_wlast,
    output wire [  USER_WIDTH-1:0] AXIM_wuser,
    output wire                    AXIM_wvalid,
    input  wire                    AXIM_wready,
    
    
    output wire [    ID_WIDTH-1:0] AXIS_bid,
    output wire [             1:0] AXIS_bresp,
    output wire [  USER_WIDTH-1:0] AXIS_buser,
    output wire                    AXIS_bvalid,
    input  wire                    AXIS_bready,
    
    input  wire [    ID_WIDTH-1:0] AXIM_bid,
    input  wire [             1:0] AXIM_bresp,
    input  wire [  USER_WIDTH-1:0] AXIM_buser,
    input  wire                    AXIM_bvalid,
    output wire                    AXIM_bready,
   
    input  wire [    ID_WIDTH-1:0] AXIS_arid,
    input  wire [  ADDR_WIDTH-1:0] AXIS_araddr,
    input  wire [   BURST_LEN-1:0] AXIS_arlen,
    input  wire [             2:0] AXIS_arsize,
    input  wire [             1:0] AXIS_arburst,
    input  wire [  LOCK_WIDTH-1:0] AXIS_arlock,
    input  wire [             3:0] AXIS_arcache,
    input  wire [             2:0] AXIS_arprot,
    input  wire [             3:0] AXIS_arregion,
    input  wire [             3:0] AXIS_arqos,
    input  wire [  USER_WIDTH-1:0] AXIS_aruser,
    input  wire                    AXIS_arvalid,
    output wire                    AXIS_arready,
   
    output wire [    ID_WIDTH-1:0] AXIM_arid,
    output wire [  ADDR_WIDTH-1:0] AXIM_araddr,
    output wire [   BURST_LEN-1:0] AXIM_arlen,
    output wire [             2:0] AXIM_arsize,
    output wire [             1:0] AXIM_arburst,
    output wire [  LOCK_WIDTH-1:0] AXIM_arlock,
    output wire [             3:0] AXIM_arcache,
    output wire [             2:0] AXIM_arprot,
    output wire [             3:0] AXIM_arregion,
    output wire [             3:0] AXIM_arqos,
    output wire [  USER_WIDTH-1:0] AXIM_aruser,
    output wire                    AXIM_arvalid,
    input  wire                    AXIM_arready,
    
    output wire [    ID_WIDTH-1:0] AXIS_rid,
    output wire [  DATA_WIDTH-1:0] AXIS_rdata,
    output wire [             1:0] AXIS_rresp,
    output wire                    AXIS_rlast,
    output wire [  USER_WIDTH-1:0] AXIS_ruser,
    output wire                    AXIS_rvalid,
    input  wire                    AXIS_rready,
    
    input  wire [    ID_WIDTH-1:0] AXIM_rid,
    input  wire [  DATA_WIDTH-1:0] AXIM_rdata,
    input  wire [             1:0] AXIM_rresp,
    input  wire                    AXIM_rlast,
    input  wire [  USER_WIDTH-1:0] AXIM_ruser,
    input  wire                    AXIM_rvalid,
    output wire                    AXIM_rready,
    // AXI stream Master (stream output wire) interface
    output wire [    ID_WIDTH-1:0] stream_tid,
    output wire [  DEST_WIDTH-1:0] stream_tdest,
    output wire [  DATA_WIDTH-1:0] stream_tdata,
    output wire [DATA_WIDTH/8-1:0] stream_tstrb,
    output wire [DATA_WIDTH/8-1:0] stream_tkeep,
    output wire                    stream_tlast,
    output wire [  USER_WIDTH-1:0] stream_tuser,
    output wire                    stream_tvalid,
    input  wire                    stream_tready
    );
    
    AXIToStream_orchestrator_Reg # (
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(ADDR_WIDTH),
      .ID_WIDTH(ID_WIDTH),
      .BURST_LEN(BURST_LEN),
      .LOCK_WIDTH(LOCK_WIDTH),
      .USER_WIDTH(USER_WIDTH),
      .DEST_WIDTH(DEST_WIDTH),
      .channels(CHANNELS)
    ) orch (
    .clk(clk),
    .resetn(resetn),
    // .RESETN_AR(RESETN_AR),
    // .RESETN_AW(RESETN_AW),
    // .RESETN_R(RESETN_R),
    // .RESETN_W(RESETN_W),
    // .RESETN_B(RESETN_B),
    .submodule_resets(submodule_resets),
    .AXIS_awid(AXIS_awid),
    .AXIS_awaddr(AXIS_awaddr),
    .AXIS_awlen(AXIS_awlen),
    .AXIS_awsize(AXIS_awsize),
    .AXIS_awburst(AXIS_awburst),
    .AXIS_awlock(AXIS_awlock),
    .AXIS_awcache(AXIS_awcache),
    .AXIS_awprot(AXIS_awprot),
    .AXIS_awregion(AXIS_awregion),
    .AXIS_awqos(AXIS_awqos),
    .AXIS_awuser(AXIS_awuser),
    .AXIS_awready(AXIS_awready),
    .AXIS_awvalid(AXIS_awvalid),
    .AXIM_awid(AXIM_awid),
    .AXIM_awaddr(AXIM_awaddr),
    .AXIM_awlen(AXIM_awlen),
    .AXIM_awsize(AXIM_awsize),
    .AXIM_awburst(AXIM_awburst),
    .AXIM_awlock(AXIM_awlock),
    .AXIM_awcache(AXIM_awcache),
    .AXIM_awprot(AXIM_awprot),
    .AXIM_awregion(AXIM_awregion),
    .AXIM_awqos(AXIM_awqos),
    .AXIM_awuser(AXIM_awuser),
    .AXIM_awready(AXIM_awready),
    .AXIM_awvalid(AXIM_awvalid),
    
    .AXIS_arid(AXIS_arid),
    .AXIS_araddr(AXIS_araddr),
    .AXIS_arlen(AXIS_arlen),
    .AXIS_arsize(AXIS_arsize),
    .AXIS_arburst(AXIS_arburst),
    .AXIS_arlock(AXIS_arlock),
    .AXIS_arcache(AXIS_arcache),
    .AXIS_arprot(AXIS_arprot),
    .AXIS_arregion(AXIS_arregion),
    .AXIS_arqos(AXIS_arqos),
    .AXIS_aruser(AXIS_aruser),
    .AXIS_arready(AXIS_arready),
    .AXIS_arvalid(AXIS_arvalid),
    .AXIM_arid(AXIM_arid),
    .AXIM_araddr(AXIM_araddr),
    .AXIM_arlen(AXIM_arlen),
    .AXIM_arsize(AXIM_arsize),
    .AXIM_arburst(AXIM_arburst),
    .AXIM_arlock(AXIM_arlock),
    .AXIM_arcache(AXIM_arcache),
    .AXIM_arprot(AXIM_arprot),
    .AXIM_arregion(AXIM_arregion),
    .AXIM_arqos(AXIM_arqos),
    .AXIM_aruser(AXIM_aruser),
    .AXIM_arready(AXIM_arready),
    .AXIM_arvalid(AXIM_arvalid),
    
    .AXIM_wid(AXIM_wid),
    .AXIM_wdata(AXIM_wdata),
    .AXIM_wstrb(AXIM_wstrb),
    .AXIM_wlast(AXIM_wlast),
    .AXIM_wuser(AXIM_wuser),
    .AXIM_wvalid(AXIM_wvalid),
    .AXIM_wready(AXIM_wready),
    .AXIS_wid(AXIS_wid),
    .AXIS_wdata(AXIS_wdata),
    .AXIS_wstrb(AXIS_wstrb),
    .AXIS_wlast(AXIS_wlast),
    .AXIS_wuser(AXIS_wuser),
    .AXIS_wvalid(AXIS_wvalid),
    .AXIS_wready(AXIS_wready),
    
    .AXIM_bid(AXIM_bid),
    .AXIM_bresp(AXIM_bresp),
    .AXIM_buser(AXIM_buser),
    .AXIM_bvalid(AXIM_bvalid),
    .AXIM_bready(AXIM_bready),
    .AXIS_bid(AXIS_bid),
    .AXIS_bresp(AXIS_bresp),
    .AXIS_buser(AXIS_buser),
    .AXIS_bvalid(AXIS_bvalid),
    .AXIS_bready(AXIS_bready),


    .AXIM_rid(AXIM_rid),
    .AXIM_rdata(AXIM_rdata),
    .AXIM_rresp(AXIM_rresp),
    .AXIM_rlast(AXIM_rlast),
    .AXIM_ruser(AXIM_ruser),
    .AXIM_rvalid(AXIM_rvalid),
    .AXIM_rready(AXIM_rready),
    .AXIS_rid(AXIS_rid),
    .AXIS_rdata(AXIS_rdata),
    .AXIS_rresp(AXIS_rresp),
    .AXIS_rlast(AXIS_rlast),
    .AXIS_ruser(AXIS_ruser),
    .AXIS_rvalid(AXIS_rvalid),
    .AXIS_rready(AXIS_rready),

    .stream_tid(stream_tid),
    .stream_tdest(stream_tdest),
    .stream_tdata(stream_tdata),
    .stream_tstrb(stream_tstrb),
    .stream_tkeep(stream_tkeep),
    .stream_tlast(stream_tlast),
    .stream_tuser(stream_tuser),
    .stream_tvalid(stream_tvalid),
    .stream_tready(stream_tready)
    );
endmodule
